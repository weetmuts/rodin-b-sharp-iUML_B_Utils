 ENTITY  Component1 IS
     port ( input_and_output_variable_declarations ) ;
 END ENTITY Component1 ;

 ARCHITECTURE Component1 IS
 	 --## <TopLevelGenerator>
 END ARCHITECTURE Component1 ;
